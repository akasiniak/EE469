module mux32to1 (out, select, muxIn);
	input logic [4:0] select;
	input logic [31:0] muxIn;
	output logic out;
	logic [1:0] outBottom4Bits;
	
	mux16to1 selectBottom4Bits1 (.out(outBottom4Bits[0]), .muxIn(muxIn[15:0]), .select(select[3:0]));
	mux16to1 selectBottom4Bits2 (.out(outBottom4Bits[1]), .muxIn(muxIn[31:16]), .select(select[3:0]));
	mux2to1 selectTopBit (.out(out), .in(outBottom4Bits), .select(select[4]));
endmodule

module mux32to1_testbench;
	logic [4:0] select;
	logic [31:0] muxIn;
	logic out;
	initial begin
		integer i;
		integer j;
		for(i = 0; i < 32; i++) begin
			select = i;
			muxIn = 1;
			for(j = 0; j < 32; j++) begin
				#10;
				muxIn = muxIn << 1;
				
			end
		end
	end
	mux32to1 dut(.out, .select, .muxIn);
endmodule